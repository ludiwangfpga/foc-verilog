`timescale 1ns / 1ps
module SimpleLogicModule (
input [15:0] a,
input [15:0] b,
input [15:0] c,
output [15:0] sum

);
reg [15:0] sin_table [0:999];
reg [15:0] cos_table [0:999];
initial begin
sin_table[0] = 16'h0000;
sin_table[1] = 16'h019C;
sin_table[2] = 16'h0337;
sin_table[3] = 16'h04D3;
sin_table[4] = 16'h066E;
sin_table[5] = 16'h0809;
sin_table[6] = 16'h09A4;
sin_table[7] = 16'h0B3F;
sin_table[8] = 16'h0CD9;
sin_table[9] = 16'h0E72;
sin_table[10] = 16'h100B;
sin_table[11] = 16'h11A3;
sin_table[12] = 16'h133A;
sin_table[13] = 16'h14D1;
sin_table[14] = 16'h1667;
sin_table[15] = 16'h17FC;
sin_table[16] = 16'h1990;
sin_table[17] = 16'h1B23;
sin_table[18] = 16'h1CB5;
sin_table[19] = 16'h1E45;
sin_table[20] = 16'h1FD5;
sin_table[21] = 16'h2163;
sin_table[22] = 16'h22F0;
sin_table[23] = 16'h247B;
sin_table[24] = 16'h2605;
sin_table[25] = 16'h278E;
sin_table[26] = 16'h2914;
sin_table[27] = 16'h2A99;
sin_table[28] = 16'h2C1D;
sin_table[29] = 16'h2D9F;
sin_table[30] = 16'h2F1E;
sin_table[31] = 16'h309C;
sin_table[32] = 16'h3218;
sin_table[33] = 16'h3392;
sin_table[34] = 16'h350A;
sin_table[35] = 16'h3680;
sin_table[36] = 16'h37F3;
sin_table[37] = 16'h3964;
sin_table[38] = 16'h3AD3;
sin_table[39] = 16'h3C40;
sin_table[40] = 16'h3DAA;
sin_table[41] = 16'h3F11;
sin_table[42] = 16'h4076;
sin_table[43] = 16'h41D9;
sin_table[44] = 16'h4338;
sin_table[45] = 16'h4495;
sin_table[46] = 16'h45F0;
sin_table[47] = 16'h4747;
sin_table[48] = 16'h489C;
sin_table[49] = 16'h49ED;
sin_table[50] = 16'h4B3C;
sin_table[51] = 16'h4C88;
sin_table[52] = 16'h4DD0;
sin_table[53] = 16'h4F15;
sin_table[54] = 16'h5058;
sin_table[55] = 16'h5196;
sin_table[56] = 16'h52D2;
sin_table[57] = 16'h540A;
sin_table[58] = 16'h553F;
sin_table[59] = 16'h5671;
sin_table[60] = 16'h579F;
sin_table[61] = 16'h58C9;
sin_table[62] = 16'h59F0;
sin_table[63] = 16'h5B13;
sin_table[64] = 16'h5C32;
sin_table[65] = 16'h5D4E;
sin_table[66] = 16'h5E66;
sin_table[67] = 16'h5F7A;
sin_table[68] = 16'h608B;
sin_table[69] = 16'h6197;
sin_table[70] = 16'h629F;
sin_table[71] = 16'h63A4;
sin_table[72] = 16'h64A4;
sin_table[73] = 16'h65A1;
sin_table[74] = 16'h6699;
sin_table[75] = 16'h678D;
sin_table[76] = 16'h687D;
sin_table[77] = 16'h6969;
sin_table[78] = 16'h6A50;
sin_table[79] = 16'h6B33;
sin_table[80] = 16'h6C12;
sin_table[81] = 16'h6CED;
sin_table[82] = 16'h6DC3;
sin_table[83] = 16'h6E94;
sin_table[84] = 16'h6F61;
sin_table[85] = 16'h702A;
sin_table[86] = 16'h70EE;
sin_table[87] = 16'h71AE;
sin_table[88] = 16'h7269;
sin_table[89] = 16'h731F;
sin_table[90] = 16'h73D0;
sin_table[91] = 16'h747D;
sin_table[92] = 16'h7526;
sin_table[93] = 16'h75C9;
sin_table[94] = 16'h7668;
sin_table[95] = 16'h7702;
sin_table[96] = 16'h7797;
sin_table[97] = 16'h7827;
sin_table[98] = 16'h78B3;
sin_table[99] = 16'h793A;
sin_table[100] = 16'h79BB;
sin_table[101] = 16'h7A38;
sin_table[102] = 16'h7AB0;
sin_table[103] = 16'h7B23;
sin_table[104] = 16'h7B91;
sin_table[105] = 16'h7BFA;
sin_table[106] = 16'h7C5D;
sin_table[107] = 16'h7CBC;
sin_table[108] = 16'h7D16;
sin_table[109] = 16'h7D6B;
sin_table[110] = 16'h7DBB;
sin_table[111] = 16'h7E05;
sin_table[112] = 16'h7E4B;
sin_table[113] = 16'h7E8B;
sin_table[114] = 16'h7EC6;
sin_table[115] = 16'h7EFD;
sin_table[116] = 16'h7F2E;
sin_table[117] = 16'h7F5A;
sin_table[118] = 16'h7F80;
sin_table[119] = 16'h7FA2;
sin_table[120] = 16'h7FBE;
sin_table[121] = 16'h7FD6;
sin_table[122] = 16'h7FE8;
sin_table[123] = 16'h7FF5;
sin_table[124] = 16'h7FFC;
sin_table[125] = 16'h7FFF;
sin_table[126] = 16'h7FFC;
sin_table[127] = 16'h7FF5;
sin_table[128] = 16'h7FE8;
sin_table[129] = 16'h7FD6;
sin_table[130] = 16'h7FBE;
sin_table[131] = 16'h7FA2;
sin_table[132] = 16'h7F80;
sin_table[133] = 16'h7F5A;
sin_table[134] = 16'h7F2E;
sin_table[135] = 16'h7EFD;
sin_table[136] = 16'h7EC6;
sin_table[137] = 16'h7E8B;
sin_table[138] = 16'h7E4B;
sin_table[139] = 16'h7E05;
sin_table[140] = 16'h7DBB;
sin_table[141] = 16'h7D6B;
sin_table[142] = 16'h7D16;
sin_table[143] = 16'h7CBC;
sin_table[144] = 16'h7C5D;
sin_table[145] = 16'h7BFA;
sin_table[146] = 16'h7B91;
sin_table[147] = 16'h7B23;
sin_table[148] = 16'h7AB0;
sin_table[149] = 16'h7A38;
sin_table[150] = 16'h79BB;
sin_table[151] = 16'h793A;
sin_table[152] = 16'h78B3;
sin_table[153] = 16'h7827;
sin_table[154] = 16'h7797;
sin_table[155] = 16'h7702;
sin_table[156] = 16'h7668;
sin_table[157] = 16'h75C9;
sin_table[158] = 16'h7526;
sin_table[159] = 16'h747D;
sin_table[160] = 16'h73D0;
sin_table[161] = 16'h731F;
sin_table[162] = 16'h7269;
sin_table[163] = 16'h71AE;
sin_table[164] = 16'h70EE;
sin_table[165] = 16'h702A;
sin_table[166] = 16'h6F61;
sin_table[167] = 16'h6E94;
sin_table[168] = 16'h6DC3;
sin_table[169] = 16'h6CED;
sin_table[170] = 16'h6C12;
sin_table[171] = 16'h6B33;
sin_table[172] = 16'h6A50;
sin_table[173] = 16'h6969;
sin_table[174] = 16'h687D;
sin_table[175] = 16'h678D;
sin_table[176] = 16'h6699;
sin_table[177] = 16'h65A1;
sin_table[178] = 16'h64A4;
sin_table[179] = 16'h63A4;
sin_table[180] = 16'h629F;
sin_table[181] = 16'h6197;
sin_table[182] = 16'h608B;
sin_table[183] = 16'h5F7A;
sin_table[184] = 16'h5E66;
sin_table[185] = 16'h5D4E;
sin_table[186] = 16'h5C32;
sin_table[187] = 16'h5B13;
sin_table[188] = 16'h59F0;
sin_table[189] = 16'h58C9;
sin_table[190] = 16'h579F;
sin_table[191] = 16'h5671;
sin_table[192] = 16'h553F;
sin_table[193] = 16'h540A;
sin_table[194] = 16'h52D2;
sin_table[195] = 16'h5196;
sin_table[196] = 16'h5058;
sin_table[197] = 16'h4F15;
sin_table[198] = 16'h4DD0;
sin_table[199] = 16'h4C88;
sin_table[200] = 16'h4B3C;
sin_table[201] = 16'h49ED;
sin_table[202] = 16'h489C;
sin_table[203] = 16'h4747;
sin_table[204] = 16'h45F0;
sin_table[205] = 16'h4495;
sin_table[206] = 16'h4338;
sin_table[207] = 16'h41D9;
sin_table[208] = 16'h4076;
sin_table[209] = 16'h3F11;
sin_table[210] = 16'h3DAA;
sin_table[211] = 16'h3C40;
sin_table[212] = 16'h3AD3;
sin_table[213] = 16'h3964;
sin_table[214] = 16'h37F3;
sin_table[215] = 16'h3680;
sin_table[216] = 16'h350A;
sin_table[217] = 16'h3392;
sin_table[218] = 16'h3218;
sin_table[219] = 16'h309C;
sin_table[220] = 16'h2F1E;
sin_table[221] = 16'h2D9F;
sin_table[222] = 16'h2C1D;
sin_table[223] = 16'h2A99;
sin_table[224] = 16'h2914;
sin_table[225] = 16'h278E;
sin_table[226] = 16'h2605;
sin_table[227] = 16'h247B;
sin_table[228] = 16'h22F0;
sin_table[229] = 16'h2163;
sin_table[230] = 16'h1FD5;
sin_table[231] = 16'h1E45;
sin_table[232] = 16'h1CB5;
sin_table[233] = 16'h1B23;
sin_table[234] = 16'h1990;
sin_table[235] = 16'h17FC;
sin_table[236] = 16'h1667;
sin_table[237] = 16'h14D1;
sin_table[238] = 16'h133A;
sin_table[239] = 16'h11A3;
sin_table[240] = 16'h100B;
sin_table[241] = 16'h0E72;
sin_table[242] = 16'h0CD9;
sin_table[243] = 16'h0B3F;
sin_table[244] = 16'h09A4;
sin_table[245] = 16'h0809;
sin_table[246] = 16'h066E;
sin_table[247] = 16'h04D3;
sin_table[248] = 16'h0337;
sin_table[249] = 16'h019C;
sin_table[250] = 16'h0000;
sin_table[251] = 16'hFE64;
sin_table[252] = 16'hFCC9;
sin_table[253] = 16'hFB2D;
sin_table[254] = 16'hF992;
sin_table[255] = 16'hF7F7;
sin_table[256] = 16'hF65C;
sin_table[257] = 16'hF4C1;
sin_table[258] = 16'hF327;
sin_table[259] = 16'hF18E;
sin_table[260] = 16'hEFF5;
sin_table[261] = 16'hEE5D;
sin_table[262] = 16'hECC6;
sin_table[263] = 16'hEB2F;
sin_table[264] = 16'hE999;
sin_table[265] = 16'hE804;
sin_table[266] = 16'hE670;
sin_table[267] = 16'hE4DD;
sin_table[268] = 16'hE34B;
sin_table[269] = 16'hE1BB;
sin_table[270] = 16'hE02B;
sin_table[271] = 16'hDE9D;
sin_table[272] = 16'hDD10;
sin_table[273] = 16'hDB85;
sin_table[274] = 16'hD9FB;
sin_table[275] = 16'hD872;
sin_table[276] = 16'hD6EC;
sin_table[277] = 16'hD567;
sin_table[278] = 16'hD3E3;
sin_table[279] = 16'hD261;
sin_table[280] = 16'hD0E2;
sin_table[281] = 16'hCF64;
sin_table[282] = 16'hCDE8;
sin_table[283] = 16'hCC6E;
sin_table[284] = 16'hCAF6;
sin_table[285] = 16'hC980;
sin_table[286] = 16'hC80D;
sin_table[287] = 16'hC69C;
sin_table[288] = 16'hC52D;
sin_table[289] = 16'hC3C0;
sin_table[290] = 16'hC256;
sin_table[291] = 16'hC0EF;
sin_table[292] = 16'hBF8A;
sin_table[293] = 16'hBE27;
sin_table[294] = 16'hBCC8;
sin_table[295] = 16'hBB6B;
sin_table[296] = 16'hBA10;
sin_table[297] = 16'hB8B9;
sin_table[298] = 16'hB764;
sin_table[299] = 16'hB613;
sin_table[300] = 16'hB4C4;
sin_table[301] = 16'hB378;
sin_table[302] = 16'hB230;
sin_table[303] = 16'hB0EB;
sin_table[304] = 16'hAFA8;
sin_table[305] = 16'hAE6A;
sin_table[306] = 16'hAD2E;
sin_table[307] = 16'hABF6;
sin_table[308] = 16'hAAC1;
sin_table[309] = 16'hA98F;
sin_table[310] = 16'hA861;
sin_table[311] = 16'hA737;
sin_table[312] = 16'hA610;
sin_table[313] = 16'hA4ED;
sin_table[314] = 16'hA3CE;
sin_table[315] = 16'hA2B2;
sin_table[316] = 16'hA19A;
sin_table[317] = 16'hA086;
sin_table[318] = 16'h9F75;
sin_table[319] = 16'h9E69;
sin_table[320] = 16'h9D61;
sin_table[321] = 16'h9C5C;
sin_table[322] = 16'h9B5C;
sin_table[323] = 16'h9A5F;
sin_table[324] = 16'h9967;
sin_table[325] = 16'h9873;
sin_table[326] = 16'h9783;
sin_table[327] = 16'h9697;
sin_table[328] = 16'h95B0;
sin_table[329] = 16'h94CD;
sin_table[330] = 16'h93EE;
sin_table[331] = 16'h9313;
sin_table[332] = 16'h923D;
sin_table[333] = 16'h916C;
sin_table[334] = 16'h909F;
sin_table[335] = 16'h8FD6;
sin_table[336] = 16'h8F12;
sin_table[337] = 16'h8E52;
sin_table[338] = 16'h8D97;
sin_table[339] = 16'h8CE1;
sin_table[340] = 16'h8C30;
sin_table[341] = 16'h8B83;
sin_table[342] = 16'h8ADA;
sin_table[343] = 16'h8A37;
sin_table[344] = 16'h8998;
sin_table[345] = 16'h88FE;
sin_table[346] = 16'h8869;
sin_table[347] = 16'h87D9;
sin_table[348] = 16'h874D;
sin_table[349] = 16'h86C6;
sin_table[350] = 16'h8645;
sin_table[351] = 16'h85C8;
sin_table[352] = 16'h8550;
sin_table[353] = 16'h84DD;
sin_table[354] = 16'h846F;
sin_table[355] = 16'h8406;
sin_table[356] = 16'h83A3;
sin_table[357] = 16'h8344;
sin_table[358] = 16'h82EA;
sin_table[359] = 16'h8295;
sin_table[360] = 16'h8245;
sin_table[361] = 16'h81FB;
sin_table[362] = 16'h81B5;
sin_table[363] = 16'h8175;
sin_table[364] = 16'h813A;
sin_table[365] = 16'h8103;
sin_table[366] = 16'h80D2;
sin_table[367] = 16'h80A6;
sin_table[368] = 16'h8080;
sin_table[369] = 16'h805E;
sin_table[370] = 16'h8042;
sin_table[371] = 16'h802A;
sin_table[372] = 16'h8018;
sin_table[373] = 16'h800B;
sin_table[374] = 16'h8004;
sin_table[375] = 16'h8001;
sin_table[376] = 16'h8004;
sin_table[377] = 16'h800B;
sin_table[378] = 16'h8018;
sin_table[379] = 16'h802A;
sin_table[380] = 16'h8042;
sin_table[381] = 16'h805E;
sin_table[382] = 16'h8080;
sin_table[383] = 16'h80A6;
sin_table[384] = 16'h80D2;
sin_table[385] = 16'h8103;
sin_table[386] = 16'h813A;
sin_table[387] = 16'h8175;
sin_table[388] = 16'h81B5;
sin_table[389] = 16'h81FB;
sin_table[390] = 16'h8245;
sin_table[391] = 16'h8295;
sin_table[392] = 16'h82EA;
sin_table[393] = 16'h8344;
sin_table[394] = 16'h83A3;
sin_table[395] = 16'h8406;
sin_table[396] = 16'h846F;
sin_table[397] = 16'h84DD;
sin_table[398] = 16'h8550;
sin_table[399] = 16'h85C8;
sin_table[400] = 16'h8645;
sin_table[401] = 16'h86C6;
sin_table[402] = 16'h874D;
sin_table[403] = 16'h87D9;
sin_table[404] = 16'h8869;
sin_table[405] = 16'h88FE;
sin_table[406] = 16'h8998;
sin_table[407] = 16'h8A37;
sin_table[408] = 16'h8ADA;
sin_table[409] = 16'h8B83;
sin_table[410] = 16'h8C30;
sin_table[411] = 16'h8CE1;
sin_table[412] = 16'h8D97;
sin_table[413] = 16'h8E52;
sin_table[414] = 16'h8F12;
sin_table[415] = 16'h8FD6;
sin_table[416] = 16'h909F;
sin_table[417] = 16'h916C;
sin_table[418] = 16'h923D;
sin_table[419] = 16'h9313;
sin_table[420] = 16'h93EE;
sin_table[421] = 16'h94CD;
sin_table[422] = 16'h95B0;
sin_table[423] = 16'h9697;
sin_table[424] = 16'h9783;
sin_table[425] = 16'h9873;
sin_table[426] = 16'h9967;
sin_table[427] = 16'h9A5F;
sin_table[428] = 16'h9B5C;
sin_table[429] = 16'h9C5C;
sin_table[430] = 16'h9D61;
sin_table[431] = 16'h9E69;
sin_table[432] = 16'h9F75;
sin_table[433] = 16'hA086;
sin_table[434] = 16'hA19A;
sin_table[435] = 16'hA2B2;
sin_table[436] = 16'hA3CE;
sin_table[437] = 16'hA4ED;
sin_table[438] = 16'hA610;
sin_table[439] = 16'hA737;
sin_table[440] = 16'hA861;
sin_table[441] = 16'hA98F;
sin_table[442] = 16'hAAC1;
sin_table[443] = 16'hABF6;
sin_table[444] = 16'hAD2E;
sin_table[445] = 16'hAE6A;
sin_table[446] = 16'hAFA8;
sin_table[447] = 16'hB0EB;
sin_table[448] = 16'hB230;
sin_table[449] = 16'hB378;
sin_table[450] = 16'hB4C4;
sin_table[451] = 16'hB613;
sin_table[452] = 16'hB764;
sin_table[453] = 16'hB8B9;
sin_table[454] = 16'hBA10;
sin_table[455] = 16'hBB6B;
sin_table[456] = 16'hBCC8;
sin_table[457] = 16'hBE27;
sin_table[458] = 16'hBF8A;
sin_table[459] = 16'hC0EF;
sin_table[460] = 16'hC256;
sin_table[461] = 16'hC3C0;
sin_table[462] = 16'hC52D;
sin_table[463] = 16'hC69C;
sin_table[464] = 16'hC80D;
sin_table[465] = 16'hC980;
sin_table[466] = 16'hCAF6;
sin_table[467] = 16'hCC6E;
sin_table[468] = 16'hCDE8;
sin_table[469] = 16'hCF64;
sin_table[470] = 16'hD0E2;
sin_table[471] = 16'hD261;
sin_table[472] = 16'hD3E3;
sin_table[473] = 16'hD567;
sin_table[474] = 16'hD6EC;
sin_table[475] = 16'hD872;
sin_table[476] = 16'hD9FB;
sin_table[477] = 16'hDB85;
sin_table[478] = 16'hDD10;
sin_table[479] = 16'hDE9D;
sin_table[480] = 16'hE02B;
sin_table[481] = 16'hE1BB;
sin_table[482] = 16'hE34B;
sin_table[483] = 16'hE4DD;
sin_table[484] = 16'hE670;
sin_table[485] = 16'hE804;
sin_table[486] = 16'hE999;
sin_table[487] = 16'hEB2F;
sin_table[488] = 16'hECC6;
sin_table[489] = 16'hEE5D;
sin_table[490] = 16'hEFF5;
sin_table[491] = 16'hF18E;
sin_table[492] = 16'hF327;
sin_table[493] = 16'hF4C1;
sin_table[494] = 16'hF65C;
sin_table[495] = 16'hF7F7;
sin_table[496] = 16'hF992;
sin_table[497] = 16'hFB2D;
sin_table[498] = 16'hFCC9;
sin_table[499] = 16'hFE64;
sin_table[500] = 16'h0000;
sin_table[501] = 16'h019C;
sin_table[502] = 16'h0337;
sin_table[503] = 16'h04D3;
sin_table[504] = 16'h066E;
sin_table[505] = 16'h0809;
sin_table[506] = 16'h09A4;
sin_table[507] = 16'h0B3F;
sin_table[508] = 16'h0CD9;
sin_table[509] = 16'h0E72;
sin_table[510] = 16'h100B;
sin_table[511] = 16'h11A3;
sin_table[512] = 16'h133A;
sin_table[513] = 16'h14D1;
sin_table[514] = 16'h1667;
sin_table[515] = 16'h17FC;
sin_table[516] = 16'h1990;
sin_table[517] = 16'h1B23;
sin_table[518] = 16'h1CB5;
sin_table[519] = 16'h1E45;
sin_table[520] = 16'h1FD5;
sin_table[521] = 16'h2163;
sin_table[522] = 16'h22F0;
sin_table[523] = 16'h247B;
sin_table[524] = 16'h2605;
sin_table[525] = 16'h278E;
sin_table[526] = 16'h2914;
sin_table[527] = 16'h2A99;
sin_table[528] = 16'h2C1D;
sin_table[529] = 16'h2D9F;
sin_table[530] = 16'h2F1E;
sin_table[531] = 16'h309C;
sin_table[532] = 16'h3218;
sin_table[533] = 16'h3392;
sin_table[534] = 16'h350A;
sin_table[535] = 16'h3680;
sin_table[536] = 16'h37F3;
sin_table[537] = 16'h3964;
sin_table[538] = 16'h3AD3;
sin_table[539] = 16'h3C40;
sin_table[540] = 16'h3DAA;
sin_table[541] = 16'h3F11;
sin_table[542] = 16'h4076;
sin_table[543] = 16'h41D9;
sin_table[544] = 16'h4338;
sin_table[545] = 16'h4495;
sin_table[546] = 16'h45F0;
sin_table[547] = 16'h4747;
sin_table[548] = 16'h489C;
sin_table[549] = 16'h49ED;
sin_table[550] = 16'h4B3C;
sin_table[551] = 16'h4C88;
sin_table[552] = 16'h4DD0;
sin_table[553] = 16'h4F15;
sin_table[554] = 16'h5058;
sin_table[555] = 16'h5196;
sin_table[556] = 16'h52D2;
sin_table[557] = 16'h540A;
sin_table[558] = 16'h553F;
sin_table[559] = 16'h5671;
sin_table[560] = 16'h579F;
sin_table[561] = 16'h58C9;
sin_table[562] = 16'h59F0;
sin_table[563] = 16'h5B13;
sin_table[564] = 16'h5C32;
sin_table[565] = 16'h5D4E;
sin_table[566] = 16'h5E66;
sin_table[567] = 16'h5F7A;
sin_table[568] = 16'h608B;
sin_table[569] = 16'h6197;
sin_table[570] = 16'h629F;
sin_table[571] = 16'h63A4;
sin_table[572] = 16'h64A4;
sin_table[573] = 16'h65A1;
sin_table[574] = 16'h6699;
sin_table[575] = 16'h678D;
sin_table[576] = 16'h687D;
sin_table[577] = 16'h6969;
sin_table[578] = 16'h6A50;
sin_table[579] = 16'h6B33;
sin_table[580] = 16'h6C12;
sin_table[581] = 16'h6CED;
sin_table[582] = 16'h6DC3;
sin_table[583] = 16'h6E94;
sin_table[584] = 16'h6F61;
sin_table[585] = 16'h702A;
sin_table[586] = 16'h70EE;
sin_table[587] = 16'h71AE;
sin_table[588] = 16'h7269;
sin_table[589] = 16'h731F;
sin_table[590] = 16'h73D0;
sin_table[591] = 16'h747D;
sin_table[592] = 16'h7526;
sin_table[593] = 16'h75C9;
sin_table[594] = 16'h7668;
sin_table[595] = 16'h7702;
sin_table[596] = 16'h7797;
sin_table[597] = 16'h7827;
sin_table[598] = 16'h78B3;
sin_table[599] = 16'h793A;
sin_table[600] = 16'h79BB;
sin_table[601] = 16'h7A38;
sin_table[602] = 16'h7AB0;
sin_table[603] = 16'h7B23;
sin_table[604] = 16'h7B91;
sin_table[605] = 16'h7BFA;
sin_table[606] = 16'h7C5D;
sin_table[607] = 16'h7CBC;
sin_table[608] = 16'h7D16;
sin_table[609] = 16'h7D6B;
sin_table[610] = 16'h7DBB;
sin_table[611] = 16'h7E05;
sin_table[612] = 16'h7E4B;
sin_table[613] = 16'h7E8B;
sin_table[614] = 16'h7EC6;
sin_table[615] = 16'h7EFD;
sin_table[616] = 16'h7F2E;
sin_table[617] = 16'h7F5A;
sin_table[618] = 16'h7F80;
sin_table[619] = 16'h7FA2;
sin_table[620] = 16'h7FBE;
sin_table[621] = 16'h7FD6;
sin_table[622] = 16'h7FE8;
sin_table[623] = 16'h7FF5;
sin_table[624] = 16'h7FFC;
sin_table[625] = 16'h7FFF;
sin_table[626] = 16'h7FFC;
sin_table[627] = 16'h7FF5;
sin_table[628] = 16'h7FE8;
sin_table[629] = 16'h7FD6;
sin_table[630] = 16'h7FBE;
sin_table[631] = 16'h7FA2;
sin_table[632] = 16'h7F80;
sin_table[633] = 16'h7F5A;
sin_table[634] = 16'h7F2E;
sin_table[635] = 16'h7EFD;
sin_table[636] = 16'h7EC6;
sin_table[637] = 16'h7E8B;
sin_table[638] = 16'h7E4B;
sin_table[639] = 16'h7E05;
sin_table[640] = 16'h7DBB;
sin_table[641] = 16'h7D6B;
sin_table[642] = 16'h7D16;
sin_table[643] = 16'h7CBC;
sin_table[644] = 16'h7C5D;
sin_table[645] = 16'h7BFA;
sin_table[646] = 16'h7B91;
sin_table[647] = 16'h7B23;
sin_table[648] = 16'h7AB0;
sin_table[649] = 16'h7A38;
sin_table[650] = 16'h79BB;
sin_table[651] = 16'h793A;
sin_table[652] = 16'h78B3;
sin_table[653] = 16'h7827;
sin_table[654] = 16'h7797;
sin_table[655] = 16'h7702;
sin_table[656] = 16'h7668;
sin_table[657] = 16'h75C9;
sin_table[658] = 16'h7526;
sin_table[659] = 16'h747D;
sin_table[660] = 16'h73D0;
sin_table[661] = 16'h731F;
sin_table[662] = 16'h7269;
sin_table[663] = 16'h71AE;
sin_table[664] = 16'h70EE;
sin_table[665] = 16'h702A;
sin_table[666] = 16'h6F61;
sin_table[667] = 16'h6E94;
sin_table[668] = 16'h6DC3;
sin_table[669] = 16'h6CED;
sin_table[670] = 16'h6C12;
sin_table[671] = 16'h6B33;
sin_table[672] = 16'h6A50;
sin_table[673] = 16'h6969;
sin_table[674] = 16'h687D;
sin_table[675] = 16'h678D;
sin_table[676] = 16'h6699;
sin_table[677] = 16'h65A1;
sin_table[678] = 16'h64A4;
sin_table[679] = 16'h63A4;
sin_table[680] = 16'h629F;
sin_table[681] = 16'h6197;
sin_table[682] = 16'h608B;
sin_table[683] = 16'h5F7A;
sin_table[684] = 16'h5E66;
sin_table[685] = 16'h5D4E;
sin_table[686] = 16'h5C32;
sin_table[687] = 16'h5B13;
sin_table[688] = 16'h59F0;
sin_table[689] = 16'h58C9;
sin_table[690] = 16'h579F;
sin_table[691] = 16'h5671;
sin_table[692] = 16'h553F;
sin_table[693] = 16'h540A;
sin_table[694] = 16'h52D2;
sin_table[695] = 16'h5196;
sin_table[696] = 16'h5058;
sin_table[697] = 16'h4F15;
sin_table[698] = 16'h4DD0;
sin_table[699] = 16'h4C88;
sin_table[700] = 16'h4B3C;
sin_table[701] = 16'h49ED;
sin_table[702] = 16'h489C;
sin_table[703] = 16'h4747;
sin_table[704] = 16'h45F0;
sin_table[705] = 16'h4495;
sin_table[706] = 16'h4338;
sin_table[707] = 16'h41D9;
sin_table[708] = 16'h4076;
sin_table[709] = 16'h3F11;
sin_table[710] = 16'h3DAA;
sin_table[711] = 16'h3C40;
sin_table[712] = 16'h3AD3;
sin_table[713] = 16'h3964;
sin_table[714] = 16'h37F3;
sin_table[715] = 16'h3680;
sin_table[716] = 16'h350A;
sin_table[717] = 16'h3392;
sin_table[718] = 16'h3218;
sin_table[719] = 16'h309C;
sin_table[720] = 16'h2F1E;
sin_table[721] = 16'h2D9F;
sin_table[722] = 16'h2C1D;
sin_table[723] = 16'h2A99;
sin_table[724] = 16'h2914;
sin_table[725] = 16'h278E;
sin_table[726] = 16'h2605;
sin_table[727] = 16'h247B;
sin_table[728] = 16'h22F0;
sin_table[729] = 16'h2163;
sin_table[730] = 16'h1FD5;
sin_table[731] = 16'h1E45;
sin_table[732] = 16'h1CB5;
sin_table[733] = 16'h1B23;
sin_table[734] = 16'h1990;
sin_table[735] = 16'h17FC;
sin_table[736] = 16'h1667;
sin_table[737] = 16'h14D1;
sin_table[738] = 16'h133A;
sin_table[739] = 16'h11A3;
sin_table[740] = 16'h100B;
sin_table[741] = 16'h0E72;
sin_table[742] = 16'h0CD9;
sin_table[743] = 16'h0B3F;
sin_table[744] = 16'h09A4;
sin_table[745] = 16'h0809;
sin_table[746] = 16'h066E;
sin_table[747] = 16'h04D3;
sin_table[748] = 16'h0337;
sin_table[749] = 16'h019C;
sin_table[750] = 16'h0000;
sin_table[751] = 16'hFE64;
sin_table[752] = 16'hFCC9;
sin_table[753] = 16'hFB2D;
sin_table[754] = 16'hF992;
sin_table[755] = 16'hF7F7;
sin_table[756] = 16'hF65C;
sin_table[757] = 16'hF4C1;
sin_table[758] = 16'hF327;
sin_table[759] = 16'hF18E;
sin_table[760] = 16'hEFF5;
sin_table[761] = 16'hEE5D;
sin_table[762] = 16'hECC6;
sin_table[763] = 16'hEB2F;
sin_table[764] = 16'hE999;
sin_table[765] = 16'hE804;
sin_table[766] = 16'hE670;
sin_table[767] = 16'hE4DD;
sin_table[768] = 16'hE34B;
sin_table[769] = 16'hE1BB;
sin_table[770] = 16'hE02B;
sin_table[771] = 16'hDE9D;
sin_table[772] = 16'hDD10;
sin_table[773] = 16'hDB85;
sin_table[774] = 16'hD9FB;
sin_table[775] = 16'hD872;
sin_table[776] = 16'hD6EC;
sin_table[777] = 16'hD567;
sin_table[778] = 16'hD3E3;
sin_table[779] = 16'hD261;
sin_table[780] = 16'hD0E2;
sin_table[781] = 16'hCF64;
sin_table[782] = 16'hCDE8;
sin_table[783] = 16'hCC6E;
sin_table[784] = 16'hCAF6;
sin_table[785] = 16'hC980;
sin_table[786] = 16'hC80D;
sin_table[787] = 16'hC69C;
sin_table[788] = 16'hC52D;
sin_table[789] = 16'hC3C0;
sin_table[790] = 16'hC256;
sin_table[791] = 16'hC0EF;
sin_table[792] = 16'hBF8A;
sin_table[793] = 16'hBE27;
sin_table[794] = 16'hBCC8;
sin_table[795] = 16'hBB6B;
sin_table[796] = 16'hBA10;
sin_table[797] = 16'hB8B9;
sin_table[798] = 16'hB764;
sin_table[799] = 16'hB613;
sin_table[800] = 16'hB4C4;
sin_table[801] = 16'hB378;
sin_table[802] = 16'hB230;
sin_table[803] = 16'hB0EB;
sin_table[804] = 16'hAFA8;
sin_table[805] = 16'hAE6A;
sin_table[806] = 16'hAD2E;
sin_table[807] = 16'hABF6;
sin_table[808] = 16'hAAC1;
sin_table[809] = 16'hA98F;
sin_table[810] = 16'hA861;
sin_table[811] = 16'hA737;
sin_table[812] = 16'hA610;
sin_table[813] = 16'hA4ED;
sin_table[814] = 16'hA3CE;
sin_table[815] = 16'hA2B2;
sin_table[816] = 16'hA19A;
sin_table[817] = 16'hA086;
sin_table[818] = 16'h9F75;
sin_table[819] = 16'h9E69;
sin_table[820] = 16'h9D61;
sin_table[821] = 16'h9C5C;
sin_table[822] = 16'h9B5C;
sin_table[823] = 16'h9A5F;
sin_table[824] = 16'h9967;
sin_table[825] = 16'h9873;
sin_table[826] = 16'h9783;
sin_table[827] = 16'h9697;
sin_table[828] = 16'h95B0;
sin_table[829] = 16'h94CD;
sin_table[830] = 16'h93EE;
sin_table[831] = 16'h9313;
sin_table[832] = 16'h923D;
sin_table[833] = 16'h916C;
sin_table[834] = 16'h909F;
sin_table[835] = 16'h8FD6;
sin_table[836] = 16'h8F12;
sin_table[837] = 16'h8E52;
sin_table[838] = 16'h8D97;
sin_table[839] = 16'h8CE1;
sin_table[840] = 16'h8C30;
sin_table[841] = 16'h8B83;
sin_table[842] = 16'h8ADA;
sin_table[843] = 16'h8A37;
sin_table[844] = 16'h8998;
sin_table[845] = 16'h88FE;
sin_table[846] = 16'h8869;
sin_table[847] = 16'h87D9;
sin_table[848] = 16'h874D;
sin_table[849] = 16'h86C6;
sin_table[850] = 16'h8645;
sin_table[851] = 16'h85C8;
sin_table[852] = 16'h8550;
sin_table[853] = 16'h84DD;
sin_table[854] = 16'h846F;
sin_table[855] = 16'h8406;
sin_table[856] = 16'h83A3;
sin_table[857] = 16'h8344;
sin_table[858] = 16'h82EA;
sin_table[859] = 16'h8295;
sin_table[860] = 16'h8245;
sin_table[861] = 16'h81FB;
sin_table[862] = 16'h81B5;
sin_table[863] = 16'h8175;
sin_table[864] = 16'h813A;
sin_table[865] = 16'h8103;
sin_table[866] = 16'h80D2;
sin_table[867] = 16'h80A6;
sin_table[868] = 16'h8080;
sin_table[869] = 16'h805E;
sin_table[870] = 16'h8042;
sin_table[871] = 16'h802A;
sin_table[872] = 16'h8018;
sin_table[873] = 16'h800B;
sin_table[874] = 16'h8004;
sin_table[875] = 16'h8001;
sin_table[876] = 16'h8004;
sin_table[877] = 16'h800B;
sin_table[878] = 16'h8018;
sin_table[879] = 16'h802A;
sin_table[880] = 16'h8042;
sin_table[881] = 16'h805E;
sin_table[882] = 16'h8080;
sin_table[883] = 16'h80A6;
sin_table[884] = 16'h80D2;
sin_table[885] = 16'h8103;
sin_table[886] = 16'h813A;
sin_table[887] = 16'h8175;
sin_table[888] = 16'h81B5;
sin_table[889] = 16'h81FB;
sin_table[890] = 16'h8245;
sin_table[891] = 16'h8295;
sin_table[892] = 16'h82EA;
sin_table[893] = 16'h8344;
sin_table[894] = 16'h83A3;
sin_table[895] = 16'h8406;
sin_table[896] = 16'h846F;
sin_table[897] = 16'h84DD;
sin_table[898] = 16'h8550;
sin_table[899] = 16'h85C8;
sin_table[900] = 16'h8645;
sin_table[901] = 16'h86C6;
sin_table[902] = 16'h874D;
sin_table[903] = 16'h87D9;
sin_table[904] = 16'h8869;
sin_table[905] = 16'h88FE;
sin_table[906] = 16'h8998;
sin_table[907] = 16'h8A37;
sin_table[908] = 16'h8ADA;
sin_table[909] = 16'h8B83;
sin_table[910] = 16'h8C30;
sin_table[911] = 16'h8CE1;
sin_table[912] = 16'h8D97;
sin_table[913] = 16'h8E52;
sin_table[914] = 16'h8F12;
sin_table[915] = 16'h8FD6;
sin_table[916] = 16'h909F;
sin_table[917] = 16'h916C;
sin_table[918] = 16'h923D;
sin_table[919] = 16'h9313;
sin_table[920] = 16'h93EE;
sin_table[921] = 16'h94CD;
sin_table[922] = 16'h95B0;
sin_table[923] = 16'h9697;
sin_table[924] = 16'h9783;
sin_table[925] = 16'h9873;
sin_table[926] = 16'h9967;
sin_table[927] = 16'h9A5F;
sin_table[928] = 16'h9B5C;
sin_table[929] = 16'h9C5C;
sin_table[930] = 16'h9D61;
sin_table[931] = 16'h9E69;
sin_table[932] = 16'h9F75;
sin_table[933] = 16'hA086;
sin_table[934] = 16'hA19A;
sin_table[935] = 16'hA2B2;
sin_table[936] = 16'hA3CE;
sin_table[937] = 16'hA4ED;
sin_table[938] = 16'hA610;
sin_table[939] = 16'hA737;
sin_table[940] = 16'hA861;
sin_table[941] = 16'hA98F;
sin_table[942] = 16'hAAC1;
sin_table[943] = 16'hABF6;
sin_table[944] = 16'hAD2E;
sin_table[945] = 16'hAE6A;
sin_table[946] = 16'hAFA8;
sin_table[947] = 16'hB0EB;
sin_table[948] = 16'hB230;
sin_table[949] = 16'hB378;
sin_table[950] = 16'hB4C4;
sin_table[951] = 16'hB613;
sin_table[952] = 16'hB764;
sin_table[953] = 16'hB8B9;
sin_table[954] = 16'hBA10;
sin_table[955] = 16'hBB6B;
sin_table[956] = 16'hBCC8;
sin_table[957] = 16'hBE27;
sin_table[958] = 16'hBF8A;
sin_table[959] = 16'hC0EF;
sin_table[960] = 16'hC256;
sin_table[961] = 16'hC3C0;
sin_table[962] = 16'hC52D;
sin_table[963] = 16'hC69C;
sin_table[964] = 16'hC80D;
sin_table[965] = 16'hC980;
sin_table[966] = 16'hCAF6;
sin_table[967] = 16'hCC6E;
sin_table[968] = 16'hCDE8;
sin_table[969] = 16'hCF64;
sin_table[970] = 16'hD0E2;
sin_table[971] = 16'hD261;
sin_table[972] = 16'hD3E3;
sin_table[973] = 16'hD567;
sin_table[974] = 16'hD6EC;
sin_table[975] = 16'hD872;
sin_table[976] = 16'hD9FB;
sin_table[977] = 16'hDB85;
sin_table[978] = 16'hDD10;
sin_table[979] = 16'hDE9D;
sin_table[980] = 16'hE02B;
sin_table[981] = 16'hE1BB;
sin_table[982] = 16'hE34B;
sin_table[983] = 16'hE4DD;
sin_table[984] = 16'hE670;
sin_table[985] = 16'hE804;
sin_table[986] = 16'hE999;
sin_table[987] = 16'hEB2F;
sin_table[988] = 16'hECC6;
sin_table[989] = 16'hEE5D;
sin_table[990] = 16'hEFF5;
sin_table[991] = 16'hF18E;
sin_table[992] = 16'hF327;
sin_table[993] = 16'hF4C1;
sin_table[994] = 16'hF65C;
sin_table[995] = 16'hF7F7;
sin_table[996] = 16'hF992;
sin_table[997] = 16'hFB2D;
sin_table[998] = 16'hFCC9;
sin_table[999] = 16'hFE64;
cos_table[0] = 16'h7FFF;
cos_table[1] = 16'h7FFC;
cos_table[2] = 16'h7FF5;
cos_table[3] = 16'h7FE8;
cos_table[4] = 16'h7FD6;
cos_table[5] = 16'h7FBE;
cos_table[6] = 16'h7FA2;
cos_table[7] = 16'h7F80;
cos_table[8] = 16'h7F5A;
cos_table[9] = 16'h7F2E;
cos_table[10] = 16'h7EFD;
cos_table[11] = 16'h7EC6;
cos_table[12] = 16'h7E8B;
cos_table[13] = 16'h7E4B;
cos_table[14] = 16'h7E05;
cos_table[15] = 16'h7DBB;
cos_table[16] = 16'h7D6B;
cos_table[17] = 16'h7D16;
cos_table[18] = 16'h7CBC;
cos_table[19] = 16'h7C5D;
cos_table[20] = 16'h7BFA;
cos_table[21] = 16'h7B91;
cos_table[22] = 16'h7B23;
cos_table[23] = 16'h7AB0;
cos_table[24] = 16'h7A38;
cos_table[25] = 16'h79BB;
cos_table[26] = 16'h793A;
cos_table[27] = 16'h78B3;
cos_table[28] = 16'h7827;
cos_table[29] = 16'h7797;
cos_table[30] = 16'h7702;
cos_table[31] = 16'h7668;
cos_table[32] = 16'h75C9;
cos_table[33] = 16'h7526;
cos_table[34] = 16'h747D;
cos_table[35] = 16'h73D0;
cos_table[36] = 16'h731F;
cos_table[37] = 16'h7269;
cos_table[38] = 16'h71AE;
cos_table[39] = 16'h70EE;
cos_table[40] = 16'h702A;
cos_table[41] = 16'h6F61;
cos_table[42] = 16'h6E94;
cos_table[43] = 16'h6DC3;
cos_table[44] = 16'h6CED;
cos_table[45] = 16'h6C12;
cos_table[46] = 16'h6B33;
cos_table[47] = 16'h6A50;
cos_table[48] = 16'h6969;
cos_table[49] = 16'h687D;
cos_table[50] = 16'h678D;
cos_table[51] = 16'h6699;
cos_table[52] = 16'h65A1;
cos_table[53] = 16'h64A4;
cos_table[54] = 16'h63A4;
cos_table[55] = 16'h629F;
cos_table[56] = 16'h6197;
cos_table[57] = 16'h608B;
cos_table[58] = 16'h5F7A;
cos_table[59] = 16'h5E66;
cos_table[60] = 16'h5D4E;
cos_table[61] = 16'h5C32;
cos_table[62] = 16'h5B13;
cos_table[63] = 16'h59F0;
cos_table[64] = 16'h58C9;
cos_table[65] = 16'h579F;
cos_table[66] = 16'h5671;
cos_table[67] = 16'h553F;
cos_table[68] = 16'h540A;
cos_table[69] = 16'h52D2;
cos_table[70] = 16'h5196;
cos_table[71] = 16'h5058;
cos_table[72] = 16'h4F15;
cos_table[73] = 16'h4DD0;
cos_table[74] = 16'h4C88;
cos_table[75] = 16'h4B3C;
cos_table[76] = 16'h49ED;
cos_table[77] = 16'h489C;
cos_table[78] = 16'h4747;
cos_table[79] = 16'h45F0;
cos_table[80] = 16'h4495;
cos_table[81] = 16'h4338;
cos_table[82] = 16'h41D9;
cos_table[83] = 16'h4076;
cos_table[84] = 16'h3F11;
cos_table[85] = 16'h3DAA;
cos_table[86] = 16'h3C40;
cos_table[87] = 16'h3AD3;
cos_table[88] = 16'h3964;
cos_table[89] = 16'h37F3;
cos_table[90] = 16'h3680;
cos_table[91] = 16'h350A;
cos_table[92] = 16'h3392;
cos_table[93] = 16'h3218;
cos_table[94] = 16'h309C;
cos_table[95] = 16'h2F1E;
cos_table[96] = 16'h2D9F;
cos_table[97] = 16'h2C1D;
cos_table[98] = 16'h2A99;
cos_table[99] = 16'h2914;
cos_table[100] = 16'h278E;
cos_table[101] = 16'h2605;
cos_table[102] = 16'h247B;
cos_table[103] = 16'h22F0;
cos_table[104] = 16'h2163;
cos_table[105] = 16'h1FD5;
cos_table[106] = 16'h1E45;
cos_table[107] = 16'h1CB5;
cos_table[108] = 16'h1B23;
cos_table[109] = 16'h1990;
cos_table[110] = 16'h17FC;
cos_table[111] = 16'h1667;
cos_table[112] = 16'h14D1;
cos_table[113] = 16'h133A;
cos_table[114] = 16'h11A3;
cos_table[115] = 16'h100B;
cos_table[116] = 16'h0E72;
cos_table[117] = 16'h0CD9;
cos_table[118] = 16'h0B3F;
cos_table[119] = 16'h09A4;
cos_table[120] = 16'h0809;
cos_table[121] = 16'h066E;
cos_table[122] = 16'h04D3;
cos_table[123] = 16'h0337;
cos_table[124] = 16'h019C;
cos_table[125] = 16'h0000;
cos_table[126] = 16'hFE64;
cos_table[127] = 16'hFCC9;
cos_table[128] = 16'hFB2D;
cos_table[129] = 16'hF992;
cos_table[130] = 16'hF7F7;
cos_table[131] = 16'hF65C;
cos_table[132] = 16'hF4C1;
cos_table[133] = 16'hF327;
cos_table[134] = 16'hF18E;
cos_table[135] = 16'hEFF5;
cos_table[136] = 16'hEE5D;
cos_table[137] = 16'hECC6;
cos_table[138] = 16'hEB2F;
cos_table[139] = 16'hE999;
cos_table[140] = 16'hE804;
cos_table[141] = 16'hE670;
cos_table[142] = 16'hE4DD;
cos_table[143] = 16'hE34B;
cos_table[144] = 16'hE1BB;
cos_table[145] = 16'hE02B;
cos_table[146] = 16'hDE9D;
cos_table[147] = 16'hDD10;
cos_table[148] = 16'hDB85;
cos_table[149] = 16'hD9FB;
cos_table[150] = 16'hD872;
cos_table[151] = 16'hD6EC;
cos_table[152] = 16'hD567;
cos_table[153] = 16'hD3E3;
cos_table[154] = 16'hD261;
cos_table[155] = 16'hD0E2;
cos_table[156] = 16'hCF64;
cos_table[157] = 16'hCDE8;
cos_table[158] = 16'hCC6E;
cos_table[159] = 16'hCAF6;
cos_table[160] = 16'hC980;
cos_table[161] = 16'hC80D;
cos_table[162] = 16'hC69C;
cos_table[163] = 16'hC52D;
cos_table[164] = 16'hC3C0;
cos_table[165] = 16'hC256;
cos_table[166] = 16'hC0EF;
cos_table[167] = 16'hBF8A;
cos_table[168] = 16'hBE27;
cos_table[169] = 16'hBCC8;
cos_table[170] = 16'hBB6B;
cos_table[171] = 16'hBA10;
cos_table[172] = 16'hB8B9;
cos_table[173] = 16'hB764;
cos_table[174] = 16'hB613;
cos_table[175] = 16'hB4C4;
cos_table[176] = 16'hB378;
cos_table[177] = 16'hB230;
cos_table[178] = 16'hB0EB;
cos_table[179] = 16'hAFA8;
cos_table[180] = 16'hAE6A;
cos_table[181] = 16'hAD2E;
cos_table[182] = 16'hABF6;
cos_table[183] = 16'hAAC1;
cos_table[184] = 16'hA98F;
cos_table[185] = 16'hA861;
cos_table[186] = 16'hA737;
cos_table[187] = 16'hA610;
cos_table[188] = 16'hA4ED;
cos_table[189] = 16'hA3CE;
cos_table[190] = 16'hA2B2;
cos_table[191] = 16'hA19A;
cos_table[192] = 16'hA086;
cos_table[193] = 16'h9F75;
cos_table[194] = 16'h9E69;
cos_table[195] = 16'h9D61;
cos_table[196] = 16'h9C5C;
cos_table[197] = 16'h9B5C;
cos_table[198] = 16'h9A5F;
cos_table[199] = 16'h9967;
cos_table[200] = 16'h9873;
cos_table[201] = 16'h9783;
cos_table[202] = 16'h9697;
cos_table[203] = 16'h95B0;
cos_table[204] = 16'h94CD;
cos_table[205] = 16'h93EE;
cos_table[206] = 16'h9313;
cos_table[207] = 16'h923D;
cos_table[208] = 16'h916C;
cos_table[209] = 16'h909F;
cos_table[210] = 16'h8FD6;
cos_table[211] = 16'h8F12;
cos_table[212] = 16'h8E52;
cos_table[213] = 16'h8D97;
cos_table[214] = 16'h8CE1;
cos_table[215] = 16'h8C30;
cos_table[216] = 16'h8B83;
cos_table[217] = 16'h8ADA;
cos_table[218] = 16'h8A37;
cos_table[219] = 16'h8998;
cos_table[220] = 16'h88FE;
cos_table[221] = 16'h8869;
cos_table[222] = 16'h87D9;
cos_table[223] = 16'h874D;
cos_table[224] = 16'h86C6;
cos_table[225] = 16'h8645;
cos_table[226] = 16'h85C8;
cos_table[227] = 16'h8550;
cos_table[228] = 16'h84DD;
cos_table[229] = 16'h846F;
cos_table[230] = 16'h8406;
cos_table[231] = 16'h83A3;
cos_table[232] = 16'h8344;
cos_table[233] = 16'h82EA;
cos_table[234] = 16'h8295;
cos_table[235] = 16'h8245;
cos_table[236] = 16'h81FB;
cos_table[237] = 16'h81B5;
cos_table[238] = 16'h8175;
cos_table[239] = 16'h813A;
cos_table[240] = 16'h8103;
cos_table[241] = 16'h80D2;
cos_table[242] = 16'h80A6;
cos_table[243] = 16'h8080;
cos_table[244] = 16'h805E;
cos_table[245] = 16'h8042;
cos_table[246] = 16'h802A;
cos_table[247] = 16'h8018;
cos_table[248] = 16'h800B;
cos_table[249] = 16'h8004;
cos_table[250] = 16'h8001;
cos_table[251] = 16'h8004;
cos_table[252] = 16'h800B;
cos_table[253] = 16'h8018;
cos_table[254] = 16'h802A;
cos_table[255] = 16'h8042;
cos_table[256] = 16'h805E;
cos_table[257] = 16'h8080;
cos_table[258] = 16'h80A6;
cos_table[259] = 16'h80D2;
cos_table[260] = 16'h8103;
cos_table[261] = 16'h813A;
cos_table[262] = 16'h8175;
cos_table[263] = 16'h81B5;
cos_table[264] = 16'h81FB;
cos_table[265] = 16'h8245;
cos_table[266] = 16'h8295;
cos_table[267] = 16'h82EA;
cos_table[268] = 16'h8344;
cos_table[269] = 16'h83A3;
cos_table[270] = 16'h8406;
cos_table[271] = 16'h846F;
cos_table[272] = 16'h84DD;
cos_table[273] = 16'h8550;
cos_table[274] = 16'h85C8;
cos_table[275] = 16'h8645;
cos_table[276] = 16'h86C6;
cos_table[277] = 16'h874D;
cos_table[278] = 16'h87D9;
cos_table[279] = 16'h8869;
cos_table[280] = 16'h88FE;
cos_table[281] = 16'h8998;
cos_table[282] = 16'h8A37;
cos_table[283] = 16'h8ADA;
cos_table[284] = 16'h8B83;
cos_table[285] = 16'h8C30;
cos_table[286] = 16'h8CE1;
cos_table[287] = 16'h8D97;
cos_table[288] = 16'h8E52;
cos_table[289] = 16'h8F12;
cos_table[290] = 16'h8FD6;
cos_table[291] = 16'h909F;
cos_table[292] = 16'h916C;
cos_table[293] = 16'h923D;
cos_table[294] = 16'h9313;
cos_table[295] = 16'h93EE;
cos_table[296] = 16'h94CD;
cos_table[297] = 16'h95B0;
cos_table[298] = 16'h9697;
cos_table[299] = 16'h9783;
cos_table[300] = 16'h9873;
cos_table[301] = 16'h9967;
cos_table[302] = 16'h9A5F;
cos_table[303] = 16'h9B5C;
cos_table[304] = 16'h9C5C;
cos_table[305] = 16'h9D61;
cos_table[306] = 16'h9E69;
cos_table[307] = 16'h9F75;
cos_table[308] = 16'hA086;
cos_table[309] = 16'hA19A;
cos_table[310] = 16'hA2B2;
cos_table[311] = 16'hA3CE;
cos_table[312] = 16'hA4ED;
cos_table[313] = 16'hA610;
cos_table[314] = 16'hA737;
cos_table[315] = 16'hA861;
cos_table[316] = 16'hA98F;
cos_table[317] = 16'hAAC1;
cos_table[318] = 16'hABF6;
cos_table[319] = 16'hAD2E;
cos_table[320] = 16'hAE6A;
cos_table[321] = 16'hAFA8;
cos_table[322] = 16'hB0EB;
cos_table[323] = 16'hB230;
cos_table[324] = 16'hB378;
cos_table[325] = 16'hB4C4;
cos_table[326] = 16'hB613;
cos_table[327] = 16'hB764;
cos_table[328] = 16'hB8B9;
cos_table[329] = 16'hBA10;
cos_table[330] = 16'hBB6B;
cos_table[331] = 16'hBCC8;
cos_table[332] = 16'hBE27;
cos_table[333] = 16'hBF8A;
cos_table[334] = 16'hC0EF;
cos_table[335] = 16'hC256;
cos_table[336] = 16'hC3C0;
cos_table[337] = 16'hC52D;
cos_table[338] = 16'hC69C;
cos_table[339] = 16'hC80D;
cos_table[340] = 16'hC980;
cos_table[341] = 16'hCAF6;
cos_table[342] = 16'hCC6E;
cos_table[343] = 16'hCDE8;
cos_table[344] = 16'hCF64;
cos_table[345] = 16'hD0E2;
cos_table[346] = 16'hD261;
cos_table[347] = 16'hD3E3;
cos_table[348] = 16'hD567;
cos_table[349] = 16'hD6EC;
cos_table[350] = 16'hD872;
cos_table[351] = 16'hD9FB;
cos_table[352] = 16'hDB85;
cos_table[353] = 16'hDD10;
cos_table[354] = 16'hDE9D;
cos_table[355] = 16'hE02B;
cos_table[356] = 16'hE1BB;
cos_table[357] = 16'hE34B;
cos_table[358] = 16'hE4DD;
cos_table[359] = 16'hE670;
cos_table[360] = 16'hE804;
cos_table[361] = 16'hE999;
cos_table[362] = 16'hEB2F;
cos_table[363] = 16'hECC6;
cos_table[364] = 16'hEE5D;
cos_table[365] = 16'hEFF5;
cos_table[366] = 16'hF18E;
cos_table[367] = 16'hF327;
cos_table[368] = 16'hF4C1;
cos_table[369] = 16'hF65C;
cos_table[370] = 16'hF7F7;
cos_table[371] = 16'hF992;
cos_table[372] = 16'hFB2D;
cos_table[373] = 16'hFCC9;
cos_table[374] = 16'hFE64;
cos_table[375] = 16'h0000;
cos_table[376] = 16'h019C;
cos_table[377] = 16'h0337;
cos_table[378] = 16'h04D3;
cos_table[379] = 16'h066E;
cos_table[380] = 16'h0809;
cos_table[381] = 16'h09A4;
cos_table[382] = 16'h0B3F;
cos_table[383] = 16'h0CD9;
cos_table[384] = 16'h0E72;
cos_table[385] = 16'h100B;
cos_table[386] = 16'h11A3;
cos_table[387] = 16'h133A;
cos_table[388] = 16'h14D1;
cos_table[389] = 16'h1667;
cos_table[390] = 16'h17FC;
cos_table[391] = 16'h1990;
cos_table[392] = 16'h1B23;
cos_table[393] = 16'h1CB5;
cos_table[394] = 16'h1E45;
cos_table[395] = 16'h1FD5;
cos_table[396] = 16'h2163;
cos_table[397] = 16'h22F0;
cos_table[398] = 16'h247B;
cos_table[399] = 16'h2605;
cos_table[400] = 16'h278E;
cos_table[401] = 16'h2914;
cos_table[402] = 16'h2A99;
cos_table[403] = 16'h2C1D;
cos_table[404] = 16'h2D9F;
cos_table[405] = 16'h2F1E;
cos_table[406] = 16'h309C;
cos_table[407] = 16'h3218;
cos_table[408] = 16'h3392;
cos_table[409] = 16'h350A;
cos_table[410] = 16'h3680;
cos_table[411] = 16'h37F3;
cos_table[412] = 16'h3964;
cos_table[413] = 16'h3AD3;
cos_table[414] = 16'h3C40;
cos_table[415] = 16'h3DAA;
cos_table[416] = 16'h3F11;
cos_table[417] = 16'h4076;
cos_table[418] = 16'h41D9;
cos_table[419] = 16'h4338;
cos_table[420] = 16'h4495;
cos_table[421] = 16'h45F0;
cos_table[422] = 16'h4747;
cos_table[423] = 16'h489C;
cos_table[424] = 16'h49ED;
cos_table[425] = 16'h4B3C;
cos_table[426] = 16'h4C88;
cos_table[427] = 16'h4DD0;
cos_table[428] = 16'h4F15;
cos_table[429] = 16'h5058;
cos_table[430] = 16'h5196;
cos_table[431] = 16'h52D2;
cos_table[432] = 16'h540A;
cos_table[433] = 16'h553F;
cos_table[434] = 16'h5671;
cos_table[435] = 16'h579F;
cos_table[436] = 16'h58C9;
cos_table[437] = 16'h59F0;
cos_table[438] = 16'h5B13;
cos_table[439] = 16'h5C32;
cos_table[440] = 16'h5D4E;
cos_table[441] = 16'h5E66;
cos_table[442] = 16'h5F7A;
cos_table[443] = 16'h608B;
cos_table[444] = 16'h6197;
cos_table[445] = 16'h629F;
cos_table[446] = 16'h63A4;
cos_table[447] = 16'h64A4;
cos_table[448] = 16'h65A1;
cos_table[449] = 16'h6699;
cos_table[450] = 16'h678D;
cos_table[451] = 16'h687D;
cos_table[452] = 16'h6969;
cos_table[453] = 16'h6A50;
cos_table[454] = 16'h6B33;
cos_table[455] = 16'h6C12;
cos_table[456] = 16'h6CED;
cos_table[457] = 16'h6DC3;
cos_table[458] = 16'h6E94;
cos_table[459] = 16'h6F61;
cos_table[460] = 16'h702A;
cos_table[461] = 16'h70EE;
cos_table[462] = 16'h71AE;
cos_table[463] = 16'h7269;
cos_table[464] = 16'h731F;
cos_table[465] = 16'h73D0;
cos_table[466] = 16'h747D;
cos_table[467] = 16'h7526;
cos_table[468] = 16'h75C9;
cos_table[469] = 16'h7668;
cos_table[470] = 16'h7702;
cos_table[471] = 16'h7797;
cos_table[472] = 16'h7827;
cos_table[473] = 16'h78B3;
cos_table[474] = 16'h793A;
cos_table[475] = 16'h79BB;
cos_table[476] = 16'h7A38;
cos_table[477] = 16'h7AB0;
cos_table[478] = 16'h7B23;
cos_table[479] = 16'h7B91;
cos_table[480] = 16'h7BFA;
cos_table[481] = 16'h7C5D;
cos_table[482] = 16'h7CBC;
cos_table[483] = 16'h7D16;
cos_table[484] = 16'h7D6B;
cos_table[485] = 16'h7DBB;
cos_table[486] = 16'h7E05;
cos_table[487] = 16'h7E4B;
cos_table[488] = 16'h7E8B;
cos_table[489] = 16'h7EC6;
cos_table[490] = 16'h7EFD;
cos_table[491] = 16'h7F2E;
cos_table[492] = 16'h7F5A;
cos_table[493] = 16'h7F80;
cos_table[494] = 16'h7FA2;
cos_table[495] = 16'h7FBE;
cos_table[496] = 16'h7FD6;
cos_table[497] = 16'h7FE8;
cos_table[498] = 16'h7FF5;
cos_table[499] = 16'h7FFC;
cos_table[500] = 16'h7FFF;
cos_table[501] = 16'h7FFC;
cos_table[502] = 16'h7FF5;
cos_table[503] = 16'h7FE8;
cos_table[504] = 16'h7FD6;
cos_table[505] = 16'h7FBE;
cos_table[506] = 16'h7FA2;
cos_table[507] = 16'h7F80;
cos_table[508] = 16'h7F5A;
cos_table[509] = 16'h7F2E;
cos_table[510] = 16'h7EFD;
cos_table[511] = 16'h7EC6;
cos_table[512] = 16'h7E8B;
cos_table[513] = 16'h7E4B;
cos_table[514] = 16'h7E05;
cos_table[515] = 16'h7DBB;
cos_table[516] = 16'h7D6B;
cos_table[517] = 16'h7D16;
cos_table[518] = 16'h7CBC;
cos_table[519] = 16'h7C5D;
cos_table[520] = 16'h7BFA;
cos_table[521] = 16'h7B91;
cos_table[522] = 16'h7B23;
cos_table[523] = 16'h7AB0;
cos_table[524] = 16'h7A38;
cos_table[525] = 16'h79BB;
cos_table[526] = 16'h793A;
cos_table[527] = 16'h78B3;
cos_table[528] = 16'h7827;
cos_table[529] = 16'h7797;
cos_table[530] = 16'h7702;
cos_table[531] = 16'h7668;
cos_table[532] = 16'h75C9;
cos_table[533] = 16'h7526;
cos_table[534] = 16'h747D;
cos_table[535] = 16'h73D0;
cos_table[536] = 16'h731F;
cos_table[537] = 16'h7269;
cos_table[538] = 16'h71AE;
cos_table[539] = 16'h70EE;
cos_table[540] = 16'h702A;
cos_table[541] = 16'h6F61;
cos_table[542] = 16'h6E94;
cos_table[543] = 16'h6DC3;
cos_table[544] = 16'h6CED;
cos_table[545] = 16'h6C12;
cos_table[546] = 16'h6B33;
cos_table[547] = 16'h6A50;
cos_table[548] = 16'h6969;
cos_table[549] = 16'h687D;
cos_table[550] = 16'h678D;
cos_table[551] = 16'h6699;
cos_table[552] = 16'h65A1;
cos_table[553] = 16'h64A4;
cos_table[554] = 16'h63A4;
cos_table[555] = 16'h629F;
cos_table[556] = 16'h6197;
cos_table[557] = 16'h608B;
cos_table[558] = 16'h5F7A;
cos_table[559] = 16'h5E66;
cos_table[560] = 16'h5D4E;
cos_table[561] = 16'h5C32;
cos_table[562] = 16'h5B13;
cos_table[563] = 16'h59F0;
cos_table[564] = 16'h58C9;
cos_table[565] = 16'h579F;
cos_table[566] = 16'h5671;
cos_table[567] = 16'h553F;
cos_table[568] = 16'h540A;
cos_table[569] = 16'h52D2;
cos_table[570] = 16'h5196;
cos_table[571] = 16'h5058;
cos_table[572] = 16'h4F15;
cos_table[573] = 16'h4DD0;
cos_table[574] = 16'h4C88;
cos_table[575] = 16'h4B3C;
cos_table[576] = 16'h49ED;
cos_table[577] = 16'h489C;
cos_table[578] = 16'h4747;
cos_table[579] = 16'h45F0;
cos_table[580] = 16'h4495;
cos_table[581] = 16'h4338;
cos_table[582] = 16'h41D9;
cos_table[583] = 16'h4076;
cos_table[584] = 16'h3F11;
cos_table[585] = 16'h3DAA;
cos_table[586] = 16'h3C40;
cos_table[587] = 16'h3AD3;
cos_table[588] = 16'h3964;
cos_table[589] = 16'h37F3;
cos_table[590] = 16'h3680;
cos_table[591] = 16'h350A;
cos_table[592] = 16'h3392;
cos_table[593] = 16'h3218;
cos_table[594] = 16'h309C;
cos_table[595] = 16'h2F1E;
cos_table[596] = 16'h2D9F;
cos_table[597] = 16'h2C1D;
cos_table[598] = 16'h2A99;
cos_table[599] = 16'h2914;
cos_table[600] = 16'h278E;
cos_table[601] = 16'h2605;
cos_table[602] = 16'h247B;
cos_table[603] = 16'h22F0;
cos_table[604] = 16'h2163;
cos_table[605] = 16'h1FD5;
cos_table[606] = 16'h1E45;
cos_table[607] = 16'h1CB5;
cos_table[608] = 16'h1B23;
cos_table[609] = 16'h1990;
cos_table[610] = 16'h17FC;
cos_table[611] = 16'h1667;
cos_table[612] = 16'h14D1;
cos_table[613] = 16'h133A;
cos_table[614] = 16'h11A3;
cos_table[615] = 16'h100B;
cos_table[616] = 16'h0E72;
cos_table[617] = 16'h0CD9;
cos_table[618] = 16'h0B3F;
cos_table[619] = 16'h09A4;
cos_table[620] = 16'h0809;
cos_table[621] = 16'h066E;
cos_table[622] = 16'h04D3;
cos_table[623] = 16'h0337;
cos_table[624] = 16'h019C;
cos_table[625] = 16'h0000;
cos_table[626] = 16'hFE64;
cos_table[627] = 16'hFCC9;
cos_table[628] = 16'hFB2D;
cos_table[629] = 16'hF992;
cos_table[630] = 16'hF7F7;
cos_table[631] = 16'hF65C;
cos_table[632] = 16'hF4C1;
cos_table[633] = 16'hF327;
cos_table[634] = 16'hF18E;
cos_table[635] = 16'hEFF5;
cos_table[636] = 16'hEE5D;
cos_table[637] = 16'hECC6;
cos_table[638] = 16'hEB2F;
cos_table[639] = 16'hE999;
cos_table[640] = 16'hE804;
cos_table[641] = 16'hE670;
cos_table[642] = 16'hE4DD;
cos_table[643] = 16'hE34B;
cos_table[644] = 16'hE1BB;
cos_table[645] = 16'hE02B;
cos_table[646] = 16'hDE9D;
cos_table[647] = 16'hDD10;
cos_table[648] = 16'hDB85;
cos_table[649] = 16'hD9FB;
cos_table[650] = 16'hD872;
cos_table[651] = 16'hD6EC;
cos_table[652] = 16'hD567;
cos_table[653] = 16'hD3E3;
cos_table[654] = 16'hD261;
cos_table[655] = 16'hD0E2;
cos_table[656] = 16'hCF64;
cos_table[657] = 16'hCDE8;
cos_table[658] = 16'hCC6E;
cos_table[659] = 16'hCAF6;
cos_table[660] = 16'hC980;
cos_table[661] = 16'hC80D;
cos_table[662] = 16'hC69C;
cos_table[663] = 16'hC52D;
cos_table[664] = 16'hC3C0;
cos_table[665] = 16'hC256;
cos_table[666] = 16'hC0EF;
cos_table[667] = 16'hBF8A;
cos_table[668] = 16'hBE27;
cos_table[669] = 16'hBCC8;
cos_table[670] = 16'hBB6B;
cos_table[671] = 16'hBA10;
cos_table[672] = 16'hB8B9;
cos_table[673] = 16'hB764;
cos_table[674] = 16'hB613;
cos_table[675] = 16'hB4C4;
cos_table[676] = 16'hB378;
cos_table[677] = 16'hB230;
cos_table[678] = 16'hB0EB;
cos_table[679] = 16'hAFA8;
cos_table[680] = 16'hAE6A;
cos_table[681] = 16'hAD2E;
cos_table[682] = 16'hABF6;
cos_table[683] = 16'hAAC1;
cos_table[684] = 16'hA98F;
cos_table[685] = 16'hA861;
cos_table[686] = 16'hA737;
cos_table[687] = 16'hA610;
cos_table[688] = 16'hA4ED;
cos_table[689] = 16'hA3CE;
cos_table[690] = 16'hA2B2;
cos_table[691] = 16'hA19A;
cos_table[692] = 16'hA086;
cos_table[693] = 16'h9F75;
cos_table[694] = 16'h9E69;
cos_table[695] = 16'h9D61;
cos_table[696] = 16'h9C5C;
cos_table[697] = 16'h9B5C;
cos_table[698] = 16'h9A5F;
cos_table[699] = 16'h9967;
cos_table[700] = 16'h9873;
cos_table[701] = 16'h9783;
cos_table[702] = 16'h9697;
cos_table[703] = 16'h95B0;
cos_table[704] = 16'h94CD;
cos_table[705] = 16'h93EE;
cos_table[706] = 16'h9313;
cos_table[707] = 16'h923D;
cos_table[708] = 16'h916C;
cos_table[709] = 16'h909F;
cos_table[710] = 16'h8FD6;
cos_table[711] = 16'h8F12;
cos_table[712] = 16'h8E52;
cos_table[713] = 16'h8D97;
cos_table[714] = 16'h8CE1;
cos_table[715] = 16'h8C30;
cos_table[716] = 16'h8B83;
cos_table[717] = 16'h8ADA;
cos_table[718] = 16'h8A37;
cos_table[719] = 16'h8998;
cos_table[720] = 16'h88FE;
cos_table[721] = 16'h8869;
cos_table[722] = 16'h87D9;
cos_table[723] = 16'h874D;
cos_table[724] = 16'h86C6;
cos_table[725] = 16'h8645;
cos_table[726] = 16'h85C8;
cos_table[727] = 16'h8550;
cos_table[728] = 16'h84DD;
cos_table[729] = 16'h846F;
cos_table[730] = 16'h8406;
cos_table[731] = 16'h83A3;
cos_table[732] = 16'h8344;
cos_table[733] = 16'h82EA;
cos_table[734] = 16'h8295;
cos_table[735] = 16'h8245;
cos_table[736] = 16'h81FB;
cos_table[737] = 16'h81B5;
cos_table[738] = 16'h8175;
cos_table[739] = 16'h813A;
cos_table[740] = 16'h8103;
cos_table[741] = 16'h80D2;
cos_table[742] = 16'h80A6;
cos_table[743] = 16'h8080;
cos_table[744] = 16'h805E;
cos_table[745] = 16'h8042;
cos_table[746] = 16'h802A;
cos_table[747] = 16'h8018;
cos_table[748] = 16'h800B;
cos_table[749] = 16'h8004;
cos_table[750] = 16'h8001;
cos_table[751] = 16'h8004;
cos_table[752] = 16'h800B;
cos_table[753] = 16'h8018;
cos_table[754] = 16'h802A;
cos_table[755] = 16'h8042;
cos_table[756] = 16'h805E;
cos_table[757] = 16'h8080;
cos_table[758] = 16'h80A6;
cos_table[759] = 16'h80D2;
cos_table[760] = 16'h8103;
cos_table[761] = 16'h813A;
cos_table[762] = 16'h8175;
cos_table[763] = 16'h81B5;
cos_table[764] = 16'h81FB;
cos_table[765] = 16'h8245;
cos_table[766] = 16'h8295;
cos_table[767] = 16'h82EA;
cos_table[768] = 16'h8344;
cos_table[769] = 16'h83A3;
cos_table[770] = 16'h8406;
cos_table[771] = 16'h846F;
cos_table[772] = 16'h84DD;
cos_table[773] = 16'h8550;
cos_table[774] = 16'h85C8;
cos_table[775] = 16'h8645;
cos_table[776] = 16'h86C6;
cos_table[777] = 16'h874D;
cos_table[778] = 16'h87D9;
cos_table[779] = 16'h8869;
cos_table[780] = 16'h88FE;
cos_table[781] = 16'h8998;
cos_table[782] = 16'h8A37;
cos_table[783] = 16'h8ADA;
cos_table[784] = 16'h8B83;
cos_table[785] = 16'h8C30;
cos_table[786] = 16'h8CE1;
cos_table[787] = 16'h8D97;
cos_table[788] = 16'h8E52;
cos_table[789] = 16'h8F12;
cos_table[790] = 16'h8FD6;
cos_table[791] = 16'h909F;
cos_table[792] = 16'h916C;
cos_table[793] = 16'h923D;
cos_table[794] = 16'h9313;
cos_table[795] = 16'h93EE;
cos_table[796] = 16'h94CD;
cos_table[797] = 16'h95B0;
cos_table[798] = 16'h9697;
cos_table[799] = 16'h9783;
cos_table[800] = 16'h9873;
cos_table[801] = 16'h9967;
cos_table[802] = 16'h9A5F;
cos_table[803] = 16'h9B5C;
cos_table[804] = 16'h9C5C;
cos_table[805] = 16'h9D61;
cos_table[806] = 16'h9E69;
cos_table[807] = 16'h9F75;
cos_table[808] = 16'hA086;
cos_table[809] = 16'hA19A;
cos_table[810] = 16'hA2B2;
cos_table[811] = 16'hA3CE;
cos_table[812] = 16'hA4ED;
cos_table[813] = 16'hA610;
cos_table[814] = 16'hA737;
cos_table[815] = 16'hA861;
cos_table[816] = 16'hA98F;
cos_table[817] = 16'hAAC1;
cos_table[818] = 16'hABF6;
cos_table[819] = 16'hAD2E;
cos_table[820] = 16'hAE6A;
cos_table[821] = 16'hAFA8;
cos_table[822] = 16'hB0EB;
cos_table[823] = 16'hB230;
cos_table[824] = 16'hB378;
cos_table[825] = 16'hB4C4;
cos_table[826] = 16'hB613;
cos_table[827] = 16'hB764;
cos_table[828] = 16'hB8B9;
cos_table[829] = 16'hBA10;
cos_table[830] = 16'hBB6B;
cos_table[831] = 16'hBCC8;
cos_table[832] = 16'hBE27;
cos_table[833] = 16'hBF8A;
cos_table[834] = 16'hC0EF;
cos_table[835] = 16'hC256;
cos_table[836] = 16'hC3C0;
cos_table[837] = 16'hC52D;
cos_table[838] = 16'hC69C;
cos_table[839] = 16'hC80D;
cos_table[840] = 16'hC980;
cos_table[841] = 16'hCAF6;
cos_table[842] = 16'hCC6E;
cos_table[843] = 16'hCDE8;
cos_table[844] = 16'hCF64;
cos_table[845] = 16'hD0E2;
cos_table[846] = 16'hD261;
cos_table[847] = 16'hD3E3;
cos_table[848] = 16'hD567;
cos_table[849] = 16'hD6EC;
cos_table[850] = 16'hD872;
cos_table[851] = 16'hD9FB;
cos_table[852] = 16'hDB85;
cos_table[853] = 16'hDD10;
cos_table[854] = 16'hDE9D;
cos_table[855] = 16'hE02B;
cos_table[856] = 16'hE1BB;
cos_table[857] = 16'hE34B;
cos_table[858] = 16'hE4DD;
cos_table[859] = 16'hE670;
cos_table[860] = 16'hE804;
cos_table[861] = 16'hE999;
cos_table[862] = 16'hEB2F;
cos_table[863] = 16'hECC6;
cos_table[864] = 16'hEE5D;
cos_table[865] = 16'hEFF5;
cos_table[866] = 16'hF18E;
cos_table[867] = 16'hF327;
cos_table[868] = 16'hF4C1;
cos_table[869] = 16'hF65C;
cos_table[870] = 16'hF7F7;
cos_table[871] = 16'hF992;
cos_table[872] = 16'hFB2D;
cos_table[873] = 16'hFCC9;
cos_table[874] = 16'hFE64;
cos_table[875] = 16'h0000;
cos_table[876] = 16'h019C;
cos_table[877] = 16'h0337;
cos_table[878] = 16'h04D3;
cos_table[879] = 16'h066E;
cos_table[880] = 16'h0809;
cos_table[881] = 16'h09A4;
cos_table[882] = 16'h0B3F;
cos_table[883] = 16'h0CD9;
cos_table[884] = 16'h0E72;
cos_table[885] = 16'h100B;
cos_table[886] = 16'h11A3;
cos_table[887] = 16'h133A;
cos_table[888] = 16'h14D1;
cos_table[889] = 16'h1667;
cos_table[890] = 16'h17FC;
cos_table[891] = 16'h1990;
cos_table[892] = 16'h1B23;
cos_table[893] = 16'h1CB5;
cos_table[894] = 16'h1E45;
cos_table[895] = 16'h1FD5;
cos_table[896] = 16'h2163;
cos_table[897] = 16'h22F0;
cos_table[898] = 16'h247B;
cos_table[899] = 16'h2605;
cos_table[900] = 16'h278E;
cos_table[901] = 16'h2914;
cos_table[902] = 16'h2A99;
cos_table[903] = 16'h2C1D;
cos_table[904] = 16'h2D9F;
cos_table[905] = 16'h2F1E;
cos_table[906] = 16'h309C;
cos_table[907] = 16'h3218;
cos_table[908] = 16'h3392;
cos_table[909] = 16'h350A;
cos_table[910] = 16'h3680;
cos_table[911] = 16'h37F3;
cos_table[912] = 16'h3964;
cos_table[913] = 16'h3AD3;
cos_table[914] = 16'h3C40;
cos_table[915] = 16'h3DAA;
cos_table[916] = 16'h3F11;
cos_table[917] = 16'h4076;
cos_table[918] = 16'h41D9;
cos_table[919] = 16'h4338;
cos_table[920] = 16'h4495;
cos_table[921] = 16'h45F0;
cos_table[922] = 16'h4747;
cos_table[923] = 16'h489C;
cos_table[924] = 16'h49ED;
cos_table[925] = 16'h4B3C;
cos_table[926] = 16'h4C88;
cos_table[927] = 16'h4DD0;
cos_table[928] = 16'h4F15;
cos_table[929] = 16'h5058;
cos_table[930] = 16'h5196;
cos_table[931] = 16'h52D2;
cos_table[932] = 16'h540A;
cos_table[933] = 16'h553F;
cos_table[934] = 16'h5671;
cos_table[935] = 16'h579F;
cos_table[936] = 16'h58C9;
cos_table[937] = 16'h59F0;
cos_table[938] = 16'h5B13;
cos_table[939] = 16'h5C32;
cos_table[940] = 16'h5D4E;
cos_table[941] = 16'h5E66;
cos_table[942] = 16'h5F7A;
cos_table[943] = 16'h608B;
cos_table[944] = 16'h6197;
cos_table[945] = 16'h629F;
cos_table[946] = 16'h63A4;
cos_table[947] = 16'h64A4;
cos_table[948] = 16'h65A1;
cos_table[949] = 16'h6699;
cos_table[950] = 16'h678D;
cos_table[951] = 16'h687D;
cos_table[952] = 16'h6969;
cos_table[953] = 16'h6A50;
cos_table[954] = 16'h6B33;
cos_table[955] = 16'h6C12;
cos_table[956] = 16'h6CED;
cos_table[957] = 16'h6DC3;
cos_table[958] = 16'h6E94;
cos_table[959] = 16'h6F61;
cos_table[960] = 16'h702A;
cos_table[961] = 16'h70EE;
cos_table[962] = 16'h71AE;
cos_table[963] = 16'h7269;
cos_table[964] = 16'h731F;
cos_table[965] = 16'h73D0;
cos_table[966] = 16'h747D;
cos_table[967] = 16'h7526;
cos_table[968] = 16'h75C9;
cos_table[969] = 16'h7668;
cos_table[970] = 16'h7702;
cos_table[971] = 16'h7797;
cos_table[972] = 16'h7827;
cos_table[973] = 16'h78B3;
cos_table[974] = 16'h793A;
cos_table[975] = 16'h79BB;
cos_table[976] = 16'h7A38;
cos_table[977] = 16'h7AB0;
cos_table[978] = 16'h7B23;
cos_table[979] = 16'h7B91;
cos_table[980] = 16'h7BFA;
cos_table[981] = 16'h7C5D;
cos_table[982] = 16'h7CBC;
cos_table[983] = 16'h7D16;
cos_table[984] = 16'h7D6B;
cos_table[985] = 16'h7DBB;
cos_table[986] = 16'h7E05;
cos_table[987] = 16'h7E4B;
cos_table[988] = 16'h7E8B;
cos_table[989] = 16'h7EC6;
cos_table[990] = 16'h7EFD;
cos_table[991] = 16'h7F2E;
cos_table[992] = 16'h7F5A;
cos_table[993] = 16'h7F80;
cos_table[994] = 16'h7FA2;
cos_table[995] = 16'h7FBE;
cos_table[996] = 16'h7FD6;
cos_table[997] = 16'h7FE8;
cos_table[998] = 16'h7FF5;
cos_table[999] = 16'h7FFC;
    end
assign sum = sin_table[a] -  cos_table[b];

endmodule
